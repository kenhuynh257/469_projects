module fetch

endmodule