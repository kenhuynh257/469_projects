module DE1_SoC(SW[0], CLOCK_50);
	input SW[0], CLOCK_50;

endmodule