module loadWord();

endmodule

module storeWord();

endmodule

module jump();

endmodule

module jumpRegister();

endmodule

module branchGreaterThan();

endmodule