module fetch ();

endmodule