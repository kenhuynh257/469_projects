module writeBack

endmodule