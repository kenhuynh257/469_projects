module hazardDetectionUnit(write_FD, write_PC, controlMux_D, memRead_DX, rs_FD, rt_FD, rt_DX);
	output write_FD, write_PC, controlMux_D;
	input memRead_DX, rs_FD, rt_FD, rt_DX;
endmodule