module instructionMemory(address,instruction);
	input[6:0] address;
	output[31:0] instruction;
	
	reg[31:0] memory[127:0];
	assign instruction = memory[address[6:0]][31:0];
	
	initial begin
	memory[0][31:0]  = 32'b000000_00000000000000000000000000; //nop
	memory[1][31:0]  = 32'b001000_01010000000000000000000011; //addi
	memory[2][31:0]  = 32'b100011_01011000000000000000000000; //lw
	memory[3][31:0]  = 32'b100011_01100000000000000000000001; //lw
	memory[4][31:0]  = 32'b100010_01111010110110000000100010; //sub
	memory[5][31:0]  = 32'b000111_01111010100000000000001101; //bgt
	memory[6][31:0]  = 32'b100011_01101000000000000000000010; //lw
	memory[7][31:0]  = 32'b000001_01101011010000000011000001; //sll
	memory[8][31:0]  = 32'b000001_01101011010000000010000001; //sll
	memory[9][31:0]  = 32'b001000_01001000000000000000000111; //addi
	memory[10][31:0] = 32'b101011_01001000000000000000000011; //sw
	memory[11][31:0] = 32'b101011_01101000000000000000000010; //sw
	memory[12][31:0] = 32'b000010_00000000000000000000010011; //j ext
	memory[13][31:0] = 32'b100011_01110000000000000000000011; //lw
	memory[14][31:0] = 32'b001000_01001000000000000000000110; //addi
	memory[15][31:0] = 32'b101011_01001000000000000000000010; //sw
	memory[16][31:0] = 32'b000001_01110011100000000010000001; //sll
	memory[17][31:0] = 32'b101011_01110000000000000000000011; //sw
	memory[18][31:0] = 32'b000010_00000000000000000000010011; //j ext
	memory[19][31:0] = 32'b000000_00000000000000000000000000; //nop ext
	memory[20][31:0] = 32'b001000_01010000000000000000000011; //addi
	memory[21][31:0] = 32'b100011_01011000000000000000000100; //lw
	memory[22][31:0] = 32'b100011_01100000000000000000000101; //lw
	memory[23][31:0] = 32'b100010_01111010110110000000100010; //sub
	memory[24][31:0] = 32'b000111_01111010100000000000100000; //bgt
	memory[25][31:0] = 32'b100011_01101000000000000000000010; //lw
	memory[26][31:0] = 32'b000001_01101011010000000011000001; //sll
	memory[27][31:0] = 32'b000001_01101011010000000010000001; //sll
	memory[28][31:0] = 32'b001000_01001000000000000000000111; //addi
	memory[29][31:0] = 32'b101011_01001000000000000000000011; //sw
	memory[30][31:0] = 32'b101011_01101000000000000000000010; //sw
	memory[31][31:0] = 32'b000010_00000000000000000000100110; //j ext2
	memory[32][31:0] = 32'b100011_01110000000000000000000011; //lw
	memory[33][31:0] = 32'b001000_01001000000000000000000110; //addi
	memory[34][31:0] = 32'b101011_01001000000000000000000010; //sw
	memory[35][31:0] = 32'b000001_01110011100000000010000001; //sll
	memory[36][31:0] = 32'b101011_01110000000000000000000011; //sw
	memory[37][31:0] = 32'b000000_00000000000000000000000000; //nop
	memory[38][31:0] = 32'b000010_00000000000000000000100110; //j ext2


	end

endmodule