module execute

endmodule