module next

endmodule