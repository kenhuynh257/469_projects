module decode ();

endmodule