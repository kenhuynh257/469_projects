module decode

endmodule